`timescale 1ms/100us

module tb_complete();

endmodule