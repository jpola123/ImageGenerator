
module image_generator (
    input logic snakeBody, snakeHead, apple, border, KeyEnc, GameOver, clk, nrst,
    output logic sync, n_cs, dc, wr, sn_rst
    output logic [7:0] D,
    output logic [3:0] x, y
);

logic [2:0] obj_code;


endmodule;